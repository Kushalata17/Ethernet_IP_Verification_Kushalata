module ab(input  a,b, output c);
  c = a+b;
endmodule
